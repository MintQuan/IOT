
module system (
	clk_clk,
	dht11_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	inout		dht11_0_external_connection_export;
	input		reset_reset_n;
endmodule
